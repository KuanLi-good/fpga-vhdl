module my_xor(in1, in2, res);
  input in1, in2;
  output res;

  assign res = in1 ^ in2;
endmodule
